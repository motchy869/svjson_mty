`ifndef JSON_PKG_DEFINED
`define JSON_PKG_DEFINED
package json_pkg;

  // Forward declarations
  typedef json_value;
  typedef json_object;
  typedef json_array;
  typedef json_string;
  typedef json_int;
  typedef json_real;
  typedef json_bool;

  // Alias to raise syntax errors in a more compact way
  `define JSON_SYNTAX_ERR(KIND, STR, IDX, DESCR="")\
    parser_result::err( \
      json_error::create( \
        .kind(KIND), \
        .description(DESCR), \
        .json_str(STR), \
        .json_pos(IDX), \
        .source_file(`__FILE__), \
        .source_line(`__LINE__) \
      ) \
    )

  // Alias to raise internal error in a more compact way
  `define JSON_INTERNAL_ERR(DESCR="", RES_T=parser_result)\
    RES_T::err( \
      json_error::create( \
        .kind(json_error::INTERNAL), \
        .description(DESCR), \
        .source_file(`__FILE__), \
        .source_line(`__LINE__) \
      ) \
    )

  // Alias to raise common error
  `define JSON_ERR(KIND, DESCR="", VAL_T=json_value)\
    json_result#(VAL_T)::err( \
      json_error::create( \
        .kind(KIND), \
        .description(DESCR), \
        .source_file(`__FILE__), \
        .source_line(`__LINE__) \
      ) \
    )

  // Utility classes
  `include "json_error.sv"
  `include "json_result.sv"

  // Interface classes for encoding standard JSON value types
  `include "encodable/json_value_encodable.sv"
  `include "encodable/json_object_encodable.sv"
  `include "encodable/json_array_encodable.sv"
  `include "encodable/json_string_encodable.sv"
  `include "encodable/json_int_encodable.sv"
  `include "encodable/json_real_encodable.sv"
  `include "encodable/json_bool_encodable.sv"

  // Wrapper classes to represent standard JSON value types
  `include "values/json_value.sv"
  `include "values/json_object.sv"
  `include "values/json_array.sv"
  `include "values/json_string.sv"
  `include "values/json_int.sv"
  `include "values/json_real.sv"
  `include "values/json_bool.sv"

  // Extension classes to handle SV specific types
  `include "values/json_enum.sv"
  `include "values/json_bits.sv"

  // JSON processors
  `include "json_decoder.sv"
  `include "json_encoder.sv"

  `undef JSON_SYNTAX_ERR
  `undef JSON_INTERNAL_ERR
  `undef JSON_ERR
endpackage : json_pkg
`endif // JSON_PKG_DEFINED
